library ieee;use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity instr_mem is
	port (
		pc1: in std_logic_vector(31 downto 0);
		pc2: in std_logic_vector(31 downto 0);
		instr1: out std_logic_vector(31 downto 0);
		instr2: out std_logic_vector(31 downto 0)
	);
end;

architecture behavior of instr_mem is
	type ramtype is array (255 downto 0) of std_logic_vector(31 downto 0);
	signal mem: ramtype;
begin

	mem(0)	<= "00100000000000010000001111111111";	--addi $1 $0 1023 
	mem(1)	<= "00111100000000100101010101010101";	--lui $2 21845    
	mem(2)	<= "00100000000000100101010101010101";	--addi $2 $0 21845
	mem(3)	<= "00111100000000110011001100110011";	--lui $3 13107    
	mem(4)	<= "00100000000000110011001100110011";	--addi $3 $0 13107
	mem(5)	<= "00111100000001000000111100001111";	--lui $4 3855     
	mem(6)	<= "00100000000001000000111100001111";	--addi $4 $0 3855
	mem(7)	<= "00000000001000000010100001000010";	--srl $5 $1 1     
	mem(8)	<= "00000000101000100010100000100100";	--and $5 $5 $2
	mem(9)	<= "00000000001001010000100000100010";	--sub $1 $1 $5
	mem(10)	<= "00000000001000110011000000100100";	--and $6 $1 $3    
	mem(11)	<= "00000000001000000011100010000010";	--srl $7 $1 2
	mem(12)	<= "00000000111000110011100000100100";	--and $7 $7 $3
	mem(13)	<= "00000000110001110000100000100000";	--add $1 $6 $7
	mem(14)	<= "00000000001000000100000100000010";	--srl $8 $1 4     
	mem(15)	<= "00000000001010000100100000100000";	--add $9 $1 $8
	mem(16)	<= "00000001001001000000100000100100";	--and $1 $9 $4
	mem(17)	<= "00000000001000000101001000000010";	--srl $10 $1 8    
	mem(18)	<= "00000000001010100000100000100000";	--add $1 $1 $10
	mem(19)	<= "00000000001000000101110000000010";	--srl $11 $1 16   
	mem(20)	<= "00000000001010110000100000100000";	--add $1 $1 $11
	mem(21)	<= "00100000000011000000000000111111";	--addi $12 $0 63  
	mem(22)	<= "00000000001011000000100000100100";	--and $1 $1 $12
	mem(23)	<= "11111111111111111111111111111111";	--exit

	process(pc1, pc2) begin
		instr1 <= mem(to_integer(unsigned(pc1(31 downto 2))));
		instr2 <= mem(to_integer(unsigned(pc2(31 downto 2))));

	end process;
end;
